`include "defines.sv"

module top(

    // Clock and Reset Inputs
    input wire clk,
    input wire rst_n,

    // Controls How Many Instructions Will be Executed
    input logic [`IMEM_ADDR_WIDTH-1:0] instruction_count
);

    // Top Level Signals
    instruction_t inst;
    wire          inst_valid;
    wire          inst_exec_begins;

    instruction_memory u_instruction_memory (
        .clk(clk),
        .rst_n(rst_n),
        .inst(inst),
        .inst_valid(inst_valid),
        .advance_pointer(inst_exec_begins),
        .instruction_count(instruction_count)
    );

    // START IMPLEMENTATION
    
    pe_inst_t pe_inst;
    wire pe_inst_valid;
    buf_inst_t buf_inst;
    wire buf_inst_valid;

    wire [`MEM0_BITWIDTH-1:0] matrix_data;
    wire [`MEM1_BITWIDTH-1:0] vector_data;
    wire [`MEM2_BITWIDTH-1:0] output_data;

    controller u_controller (
        .clk(clk),
    .rst_n(rst_n),

    .inst(inst),
    .inst_valid(inst_valid),
    .inst_exec_begins(inst_exec_begins),

    .pe_inst(pe_inst),
    .pe_inst_valid(pe_inst_valid),
    .buf_inst(buf_inst),
    .buf_inst_valid(buf_inst_valid)
    );

    buffer u_buffer (
        .clk(clk),
    .rst_n(rst_n),

    .buf_inst(buf_inst),
    .buf_inst_valid(buf_inst_valid),

    .matrix_data(matrix_data),
    .vector_data(vector_data),
    .output_data(output_data)
    );

    wire [`PE_OUTPUT_BITWIDTH-1:0] vector_output [`PE_COUNT-1:0];

    genvar i;

    generate
        for (i = 0; i < `PE_COUNT; i = i + 1) begin  
                  processing_element u_processing_element ( 
                      .clk(clk),
                      .rst_n(rst_n),
                      .pe_inst(pe_inst),
                      .pe_inst_valid(pe_inst_valid),
                          .vector_input(vector_data),
                          .matrix_input(matrix_data[`MEM0_BITWIDTH-1 - i*`PE_INPUT_BITWIDTH -: `PE_INPUT_BITWIDTH]),
                          .vector_output(vector_output[i])
              );
        end
    endgenerate

    genvar j;
    generate
      for (j = 0; j < `PE_COUNT; j = j + 1) begin 
        assign output_data[`MEM2_BITWIDTH-1 - j*`PE_OUTPUT_BITWIDTH -: `PE_OUTPUT_BITWIDTH] = vector_output[j];

   end
   endgenerate  
    // END IMPLEMENTATION
endmodule

